module Adder_2
(
    input [63:0] A, B,
    output [63:0] out
);

assign out = A + B;

endmodule // Adder
